.model xxxxxxxx D
+ IS=2.939E-13
+ N=4.0113
+ RS=0.24229
+ EG=3
+ XIT=25
*$